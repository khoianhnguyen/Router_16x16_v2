`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/30/2024 01:42:04 PM
// Design Name: 
// Module Name: router
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module router
   (clk,
    din,
    frame_n,
    reset_n,
    valid_n,
    frame_o,
    valid_o,
    dout);
  input clk;
  input [15:0]din;
  input [15:0]frame_n;
  input [15:0] valid_n;
  output [15:0] frame_o;
  output [15:0] valid_o;
  output [15:0] dout; 
  input reset_n;
  wire clk_1;
  wire [15:0]matrix_0_dout0;
  wire [15:0]matrix_0_dout1;
  wire [15:0]matrix_0_dout10;
  wire [15:0]matrix_0_dout11;
  wire [15:0]matrix_0_dout12;
  wire [15:0]matrix_0_dout13;
  wire [15:0]matrix_0_dout14;
  wire [15:0]matrix_0_dout15;
  wire [15:0]matrix_0_dout2;
  wire [15:0]matrix_0_dout3;
  wire [15:0]matrix_0_dout4;
  wire [15:0]matrix_0_dout5;
  wire [15:0]matrix_0_dout6;
  wire [15:0]matrix_0_dout7;
  wire [15:0]matrix_0_dout8;
  wire [15:0]matrix_0_dout9;
  wire [15:0]matrix_0_frame_o0;
  wire [15:0]matrix_0_frame_o1;
  wire [15:0]matrix_0_frame_o10;
  wire [15:0]matrix_0_frame_o11;
  wire [15:0]matrix_0_frame_o12;
  wire [15:0]matrix_0_frame_o13;
  wire [15:0]matrix_0_frame_o14;
  wire [15:0]matrix_0_frame_o15;
  wire [15:0]matrix_0_frame_o2;
  wire [15:0]matrix_0_frame_o3;
  wire [15:0]matrix_0_frame_o4;
  wire [15:0]matrix_0_frame_o5;
  wire [15:0]matrix_0_frame_o6;
  wire [15:0]matrix_0_frame_o7;
  wire [15:0]matrix_0_frame_o8;
  wire [15:0]matrix_0_frame_o9;
  wire [15:0]matrix_0_request_o0;
  wire [15:0]matrix_0_request_o1;
  wire [15:0]matrix_0_request_o10;
  wire [15:0]matrix_0_request_o11;
  wire [15:0]matrix_0_request_o12;
  wire [15:0]matrix_0_request_o13;
  wire [15:0]matrix_0_request_o14;
  wire [15:0]matrix_0_request_o15;
  wire [15:0]matrix_0_request_o2;
  wire [15:0]matrix_0_request_o3;
  wire [15:0]matrix_0_request_o4;
  wire [15:0]matrix_0_request_o5;
  wire [15:0]matrix_0_request_o6;
  wire [15:0]matrix_0_request_o7;
  wire [15:0]matrix_0_request_o8;
  wire [15:0]matrix_0_request_o9;
  wire [15:0]matrix_0_valid_o0;
  wire [15:0]matrix_0_valid_o1;
  wire [15:0]matrix_0_valid_o10;
  wire [15:0]matrix_0_valid_o11;
  wire [15:0]matrix_0_valid_o12;
  wire [15:0]matrix_0_valid_o13;
  wire [15:0]matrix_0_valid_o14;
  wire [15:0]matrix_0_valid_o15;
  wire [15:0]matrix_0_valid_o2;
  wire [15:0]matrix_0_valid_o3;
  wire [15:0]matrix_0_valid_o4;
  wire [15:0]matrix_0_valid_o5;
  wire [15:0]matrix_0_valid_o6;
  wire [15:0]matrix_0_valid_o7;
  wire [15:0]matrix_0_valid_o8;
  wire [15:0]matrix_0_valid_o9;
  wire reset_n_1;
  wire [15:0]router2decode_0_dout;
  wire [15:0]router2decode_0_frame_o;
  wire [15:0]router2decode_0_request;
  wire [15:0]router2decode_0_valid_o;
  wire [15:0]router2decode_10_dout;
  wire [15:0]router2decode_10_frame_o;
  wire [15:0]router2decode_10_request;
  wire [15:0]router2decode_10_valid_o;
  wire [15:0]router2decode_11_dout;
  wire [15:0]router2decode_11_frame_o;
  wire [15:0]router2decode_11_request;
  wire [15:0]router2decode_11_valid_o;
  wire [15:0]router2decode_12_dout;
  wire [15:0]router2decode_12_frame_o;
  wire [15:0]router2decode_12_request;
  wire [15:0]router2decode_12_valid_o;
  wire [15:0]router2decode_13_dout;
  wire [15:0]router2decode_13_frame_o;
  wire [15:0]router2decode_13_request;
  wire [15:0]router2decode_13_valid_o;
  wire [15:0]router2decode_14_dout;
  wire [15:0]router2decode_14_frame_o;
  wire [15:0]router2decode_14_request;
  wire [15:0]router2decode_14_valid_o;
  wire [15:0]router2decode_15_dout;
  wire [15:0]router2decode_15_frame_o;
  wire [15:0]router2decode_15_request;
  wire [15:0]router2decode_15_valid_o;
  wire [15:0]router2decode_1_dout;
  wire [15:0]router2decode_1_frame_o;
  wire [15:0]router2decode_1_request;
  wire [15:0]router2decode_1_valid_o;
  wire [15:0]router2decode_2_dout;
  wire [15:0]router2decode_2_frame_o;
  wire [15:0]router2decode_2_request;
  wire [15:0]router2decode_2_valid_o;
  wire [15:0]router2decode_3_dout;
  wire [15:0]router2decode_3_frame_o;
  wire [15:0]router2decode_3_request;
  wire [15:0]router2decode_3_valid_o;
  wire [15:0]router2decode_4_dout;
  wire [15:0]router2decode_4_frame_o;
  wire [15:0]router2decode_4_request;
  wire [15:0]router2decode_4_valid_o;
  wire [15:0]router2decode_5_dout;
  wire [15:0]router2decode_5_frame_o;
  wire [15:0]router2decode_5_request;
  wire [15:0]router2decode_5_valid_o;
  wire [15:0]router2decode_6_dout;
  wire [15:0]router2decode_6_frame_o;
  wire [15:0]router2decode_6_request;
  wire [15:0]router2decode_6_valid_o;
  wire [15:0]router2decode_7_dout;
  wire [15:0]router2decode_7_frame_o;
  wire [15:0]router2decode_7_request;
  wire [15:0]router2decode_7_valid_o;
  wire [15:0]router2decode_8_dout;
  wire [15:0]router2decode_8_frame_o;
  wire [15:0]router2decode_8_request;
  wire [15:0]router2decode_8_valid_o;
  wire [15:0]router2decode_9_dout;
  wire [15:0]router2decode_9_frame_o;
  wire [15:0]router2decode_9_request;
  wire [15:0]router2decode_9_valid_o;

  assign clk_1 = clk;
  assign reset_n_1 = reset_n;
  arbiter2enable_wrapper arbiter2enable_wrapp_0
       (.din(matrix_0_dout0),
        .frame_n(matrix_0_frame_o0),
        .request(matrix_0_request_o0),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o0),
        .dout(dout[0]),
        .frame_o(frame_o[0]),
        .valid_o(valid_o[0]));
  arbiter2enable_wrapper arbiter2enable_wrapp_1
       (.din(matrix_0_dout1),
        .frame_n(matrix_0_frame_o1),
        .request(matrix_0_request_o1),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o1),
        .dout(dout[1]),
        .frame_o(frame_o[1]),
        .valid_o(valid_o[1]));
  arbiter2enable_wrapper arbiter2enable_wrapp_2
       (.din(matrix_0_dout2),
        .frame_n(matrix_0_frame_o2),
        .request(matrix_0_request_o2),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o2),
        .dout(dout[2]),
        .frame_o(frame_o[2]),
        .valid_o(valid_o[2]));
  arbiter2enable_wrapper arbiter2enable_wrapp_3
       (.din(matrix_0_dout3),
        .frame_n(matrix_0_frame_o3),
        .request(matrix_0_request_o3),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o3),
        .dout(dout[3]),
        .frame_o(frame_o[3]),
        .valid_o(valid_o[3]));
  arbiter2enable_wrapper arbiter2enable_wrapp_4
       (.din(matrix_0_dout4),
        .frame_n(matrix_0_frame_o4),
        .request(matrix_0_request_o4),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o4),
        .dout(dout[4]),
        .frame_o(frame_o[4]),
        .valid_o(valid_o[4]));
  arbiter2enable_wrapper arbiter2enable_wrapp_5
       (.din(matrix_0_dout5),
        .frame_n(matrix_0_frame_o5),
        .request(matrix_0_request_o5),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o5),
        .dout(dout[5]),
        .frame_o(frame_o[5]),
        .valid_o(valid_o[5]));
  arbiter2enable_wrapper arbiter2enable_wrapp_6
       (.din(matrix_0_dout6),
        .frame_n(matrix_0_frame_o6),
        .request(matrix_0_request_o6),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o6),
        .dout(dout[6]),
        .frame_o(frame_o[6]),
        .valid_o(valid_o[6]));
  arbiter2enable_wrapper arbiter2enable_wrapp_7
       (.din(matrix_0_dout7),
        .frame_n(matrix_0_frame_o7),
        .request(matrix_0_request_o7),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o7),
        .dout(dout[7]),
        .frame_o(frame_o[7]),
        .valid_o(valid_o[7]));
  arbiter2enable_wrapper arbiter2enable_wrapp_8
       (.din(matrix_0_dout8),
        .frame_n(matrix_0_frame_o8),
        .request(matrix_0_request_o8),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o8),
        .dout(dout[8]),
        .frame_o(frame_o[8]),
        .valid_o(valid_o[8]));
  arbiter2enable_wrapper arbiter2enable_wrapp_9
       (.din(matrix_0_dout2),
        .frame_n(matrix_0_frame_o9),
        .request(matrix_0_request_o9),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o9),
        .dout(dout[9]),
        .frame_o(frame_o[9]),
        .valid_o(valid_o[9]));
  arbiter2enable_wrapper arbiter2enable_wrapp_10
       (.din(matrix_0_dout10),
        .frame_n(matrix_0_frame_o10),
        .request(matrix_0_request_o10),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o10),
        .dout(dout[10]),
        .frame_o(frame_o[10]),
        .valid_o(valid_o[10]));
  arbiter2enable_wrapper arbiter2enable_wrapp_11
       (.din(matrix_0_dout11),
        .frame_n(matrix_0_frame_o11),
        .request(matrix_0_request_o11),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o11),
        .dout(dout[11]),
        .frame_o(frame_o[11]),
        .valid_o(valid_o[11]));
  arbiter2enable_wrapper arbiter2enable_wrapp_12
       (.din(matrix_0_dout12),
        .frame_n(matrix_0_frame_o12),
        .request(matrix_0_request_o12),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o12),
        .dout(dout[12]),
        .frame_o(frame_o[12]),
        .valid_o(valid_o[12]));
  arbiter2enable_wrapper arbiter2enable_wrapp_13
       (.din(matrix_0_dout13),
        .frame_n(matrix_0_frame_o13),
        .request(matrix_0_request_o13),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o13),
        .dout(dout[13]),
        .frame_o(frame_o[13]),
        .valid_o(valid_o[13]));
  arbiter2enable_wrapper arbiter2enable_wrapp_14
       (.din(matrix_0_dout14),
        .frame_n(matrix_0_frame_o14),
        .request(matrix_0_request_o14),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o14),
        .dout(dout[14]),
        .frame_o(frame_o[14]),
        .valid_o(valid_o[14]));
  arbiter2enable_wrapper arbiter2enable_wrapp_15
       (.din(matrix_0_dout15),
        .frame_n(matrix_0_frame_15),
        .request(matrix_0_request_o15),
        .reset_n(reset_n_1),
        .valid_n(matrix_0_valid_o15),
        .dout(dout[15]),
        .frame_o(frame_o[15]),
        .valid_o(valid_o[15]));
  matrix matrix_0
       (.din0(router2decode_0_dout),
        .din1(router2decode_1_dout),
        .din10(router2decode_10_dout),
        .din11(router2decode_11_dout),
        .din12(router2decode_12_dout),
        .din13(router2decode_12_dout),
        .din14(router2decode_14_dout),
        .din15(router2decode_15_dout),
        .din2(router2decode_2_dout),
        .din3(router2decode_3_dout),
        .din4(router2decode_4_dout),
        .din5(router2decode_5_dout),
        .din6(router2decode_6_dout),
        .din7(router2decode_7_dout),
        .din8(router2decode_8_dout),
        .din9(router2decode_9_dout),
        .dout0(matrix_0_dout0),
        .dout1(matrix_0_dout1),
        .dout10(matrix_0_dout10),
        .dout11(matrix_0_dout11),
        .dout12(matrix_0_dout12),
        .dout13(matrix_0_dout13),
        .dout14(matrix_0_dout14),
        .dout15(matrix_0_dout15),
        .dout2(matrix_0_dout2),
        .dout3(matrix_0_dout3),
        .dout4(matrix_0_dout4),
        .dout5(matrix_0_dout5),
        .dout6(matrix_0_dout6),
        .dout7(matrix_0_dout7),
        .dout8(matrix_0_dout8),
        .dout9(matrix_0_dout9),
        .frame_n0(router2decode_0_frame_o),
        .frame_n1(router2decode_1_frame_o),
        .frame_n10(router2decode_10_frame_o),
        .frame_n11(router2decode_11_frame_o),
        .frame_n12(router2decode_12_frame_o),
        .frame_n13(router2decode_13_frame_o),
        .frame_n14(router2decode_14_frame_o),
        .frame_n15(router2decode_15_frame_o),
        .frame_n2(router2decode_2_frame_o),
        .frame_n3(router2decode_3_frame_o),
        .frame_n4(router2decode_4_frame_o),
        .frame_n5(router2decode_5_frame_o),
        .frame_n6(router2decode_6_frame_o),
        .frame_n7(router2decode_7_frame_o),
        .frame_n8(router2decode_8_frame_o),
        .frame_n9(router2decode_9_frame_o),
        .frame_o0(matrix_0_frame_o0),
        .frame_o1(matrix_0_frame_o1),
        .frame_o10(matrix_0_frame_o10),
        .frame_o11(matrix_0_frame_o11),
        .frame_o12(matrix_0_frame_o12),
        .frame_o13(matrix_0_frame_o13),
        .frame_o14(matrix_0_frame_o14),
        .frame_o15(matrix_0_frame_o15),
        .frame_o2(matrix_0_frame_o2),
        .frame_o3(matrix_0_frame_o3),
        .frame_o4(matrix_0_frame_o4),
        .frame_o5(matrix_0_frame_o5),
        .frame_o6(matrix_0_frame_o6),
        .frame_o7(matrix_0_frame_o7),
        .frame_o8(matrix_0_frame_o8),
        .frame_o9(matrix_0_frame_o9),
        .request0(router2decode_0_request),
        .request1(router2decode_1_request),
        .request10(router2decode_10_request),
        .request11(router2decode_11_request),
        .request12(router2decode_12_request),
        .request13(router2decode_13_request),
        .request14(router2decode_14_request),
        .request15(router2decode_15_request),
        .request2(router2decode_2_request),
        .request3(router2decode_3_request),
        .request4(router2decode_4_request),
        .request5(router2decode_5_request),
        .request6(router2decode_6_request),
        .request7(router2decode_7_request),
        .request8(router2decode_8_request),
        .request9(router2decode_9_request),
        .request_o0(matrix_0_request_o0),
        .request_o1(matrix_0_request_o1),
        .request_o10(matrix_0_request_o10),
        .request_o11(matrix_0_request_o11),
        .request_o12(matrix_0_request_o12),
        .request_o13(matrix_0_request_o13),
        .request_o14(matrix_0_request_o14),
        .request_o15(matrix_0_request_o15),
        .request_o2(matrix_0_request_o2),
        .request_o3(matrix_0_request_o3),
        .request_o4(matrix_0_request_o4),
        .request_o5(matrix_0_request_o5),
        .request_o6(matrix_0_request_o6),
        .request_o7(matrix_0_request_o7),
        .request_o8(matrix_0_request_o8),
        .request_o9(matrix_0_request_o9),
        .valid_n0(router2decode_0_valid_o),
        .valid_n1(router2decode_1_valid_o),
        .valid_n10(router2decode_10_valid_o),
        .valid_n11(router2decode_11_valid_o),
        .valid_n12(router2decode_12_valid_o),
        .valid_n13(router2decode_13_valid_o),
        .valid_n14(router2decode_14_valid_o),
        .valid_n15(router2decode_15_valid_o),
        .valid_n2(router2decode_2_valid_o),
        .valid_n3(router2decode_3_valid_o),
        .valid_n4(router2decode_4_valid_o),
        .valid_n5(router2decode_5_valid_o),
        .valid_n6(router2decode_6_valid_o),
        .valid_n7(router2decode_7_valid_o),
        .valid_n8(router2decode_8_valid_o),
        .valid_n9(router2decode_9_valid_o),
        .valid_o0(matrix_0_valid_o0),
        .valid_o1(matrix_0_valid_o1),
        .valid_o10(matrix_0_valid_o10),
        .valid_o11(matrix_0_valid_o11),
        .valid_o12(matrix_0_valid_o12),
        .valid_o13(matrix_0_valid_o13),
        .valid_o14(matrix_0_valid_o14),
        .valid_o15(matrix_0_valid_o15),
        .valid_o2(matrix_0_valid_o2),
        .valid_o3(matrix_0_valid_o3),
        .valid_o4(matrix_0_valid_o4),
        .valid_o5(matrix_0_valid_o5),
        .valid_o6(matrix_0_valid_o6),
        .valid_o7(matrix_0_valid_o7),
        .valid_o8(matrix_0_valid_o8),
        .valid_o9(matrix_0_valid_o9));
  router2decode router2decode_0
       (.clk(clk_1),
        .din(din[0]),
        .dout(router2decode_0_dout),
        .frame_n(frame_n[0]),
        .frame_o(router2decode_0_frame_o),
        .request(router2decode_0_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[0]),
        .valid_o(router2decode_0_valid_o));
  router2decode router2decode_1
       (.clk(clk_1),
        .din(din[1]),
        .dout(router2decode_1_dout),
        .frame_n(frame_n[1]),
        .frame_o(router2decode_1_frame_o),
        .request(router2decode_1_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[1]),
        .valid_o(router2decode_1_valid_o));
  router2decode router2decode_2
       (.clk(clk_1),
        .din(din[2]),
        .dout(router2decode_2_dout),
        .frame_n(frame_n[2]),
        .frame_o(router2decode_2_frame_o),
        .request(router2decode_2_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[2]),
        .valid_o(router2decode_2_valid_o));
  router2decode router2decode_3
       (.clk(clk_1),
        .din(din[3]),
        .dout(router2decode_3_dout),
        .frame_n(frame_n[3]),
        .frame_o(router2decode_3_frame_o),
        .request(router2decode_3_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[3]),
        .valid_o(router2decode_3_valid_o));
  router2decode router2decode_4
       (.clk(clk_1),
        .din(din[4]),
        .dout(router2decode_4_dout),
        .frame_n(frame_n[4]),
        .frame_o(router2decode_4_frame_o),
        .request(router2decode_4_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[4]),
        .valid_o(router2decode_4_valid_o));
  router2decode router2decode_5
       (.clk(clk_1),
        .din(din[5]),
        .dout(router2decode_5_dout),
        .frame_n(frame_n[5]),
        .frame_o(router2decode_5_frame_o),
        .request(router2decode_5_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[5]),
        .valid_o(router2decode_5_valid_o));
  router2decode router2decode_6
       (.clk(clk_1),
        .din(din[6]),
        .dout(router2decode_6_dout),
        .frame_n(frame_n[6]),
        .frame_o(router2decode_6_frame_o),
        .request(router2decode_6_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[6]),
        .valid_o(router2decode_6_valid_o));
  router2decode router2decode_7
       (.clk(clk_1),
        .din(din[7]),
        .dout(router2decode_7_dout),
        .frame_n(frame_n[7]),
        .frame_o(router2decode_7_frame_o),
        .request(router2decode_7_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[7]),
        .valid_o(router2decode_7_valid_o));
  router2decode router2decode_8
       (.clk(clk_1),
        .din(din[8]),
        .dout(router2decode_8_dout),
        .frame_n(frame_n[8]),
        .frame_o(router2decode_8_frame_o),
        .request(router2decode_8_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[8]),
        .valid_o(router2decode_8_valid_o));
  router2decode router2decode_9
       (.clk(clk_1),
        .din(din[9]),
        .dout(router2decode_9_dout),
        .frame_n(frame_n[9]),
        .frame_o(router2decode_9_frame_o),
        .request(router2decode_9_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[9]),
        .valid_o(router2decode_9_valid_o));
  router2decode router2decode_10
       (.clk(clk_1),
        .din(din[10]),
        .dout(router2decode_10_dout),
        .frame_n(frame_n[10]),
        .frame_o(router2decode_10_frame_o),
        .request(router2decode_10_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[10]),
        .valid_o(router2decode_10_valid_o));
  router2decode router2decode_11
       (.clk(clk_1),
        .din(din[11]),
        .dout(router2decode_11_dout),
        .frame_n(frame_n[11]),
        .frame_o(router2decode_11_frame_o),
        .request(router2decode_11_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[11]),
        .valid_o(router2decode_11_valid_o));
  router2decode router2decode_12
       (.clk(clk_1),
        .din(din[12]),
        .dout(router2decode_12_dout),
        .frame_n(frame_n[12]),
        .frame_o(router2decode_12_frame_o),
        .request(router2decode_12_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[12]),
        .valid_o(router2decode_12_valid_o));
  router2decode router2decode_13
       (.clk(clk_1),
        .din(din[13]),
        .dout(router2decode_13_dout),
        .frame_n(frame_n[13]),
        .frame_o(router2decode_13_frame_o),
        .request(router2decode_13_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[13]),
        .valid_o(router2decode_13_valid_o));
  router2decode router2decode_14
       (.clk(clk_1),
        .din(din[14]),
        .dout(router2decode_14_dout),
        .frame_n(frame_n[14]),
        .frame_o(router2decode_14_frame_o),
        .request(router2decode_14_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[14]),
        .valid_o(router2decode_14_valid_o));
  router2decode router2decode_15
       (.clk(clk_1),
        .din(din[15]),
        .dout(router2decode_15_dout),
        .frame_n(frame_n[15]),
        .frame_o(router2decode_15_frame_o),
        .request(router2decode_15_request),
        .reset_n(reset_n_1),
        .valid_n(valid_n[15]),
        .valid_o(router2decode_15_valid_o));
endmodule
